`ifndef CONFIGURATION_PKG_SV
`define CONFIGURATION_PKG_SV

package configurations_pkg;

   import uvm_pkg::*;      // import the UVM library   
 `include "uvm_macros.svh" // Include the UVM macros

`include "file_cnn_config.sv"


endpackage : configurations_pkg

`endif
